`define OPCODE_BRANCH 7'b1100011

module IFetch(
    input wire clk,
    input wire rst,
    input wire rdy,

    input wire rollback
)

endmodule