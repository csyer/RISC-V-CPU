module ROB(
    input wire clk,
    input wire rst,
    input wire rdy
);

always @(posedge clk) begin
    if (rst) begin
        // TODO
    end else if (rdy) begin
        // TODO
    end
end

endmodule