// RISCV32I CPU top module
// port modification allowed for debugging purposes

`include "memctrl.v"

module cpu(
    input  wire                 clk_in,			// system clock signal
    input  wire                 rst_in,			// reset signal
	input  wire					        rdy_in,			// ready signal, pause cpu when low

    input  wire [ 7:0]          mem_din,		// data input bus
    output wire [ 7:0]          mem_dout,		// data output bus
    output wire [31:0]          mem_a,			// address bus (only 17:0 is used)
    output wire                 mem_wr,			// write/read signal (1 for write)
	
	input  wire                 io_buffer_full, // 1 if uart buffer is full
	
	output wire [31:0]			dbgreg_dout		// cpu register output (debugging demo)
);

// implementation goes here

// Specifications:
// - Pause cpu(freeze pc, registers, etc.) when rdy_in is low
// - Memory read result will be returned in the next cycle. Write takes 1 cycle(no need to wait)
// - Memory is of size 128KB, with valid address ranging from 0x0 to 0x20000
// - I/O port is mapped to address higher than 0x30000 (mem_a[17:16]==2'b11)
// - 0x30000 read: read a byte from input
// - 0x30000 write: write a byte to output (write 0x00 is ignored)
// - 0x30004 read: read clocks passed since cpu starts (in dword, 4 bytes)
// - 0x30004 write: indicates program stop (will output '\0' through uart tx)

wire rollback;

wire if_to_mem_en;
wire [`ADDR_WID] if_to_mem_pc;
wire mem_to_if_done;
wire [`ICACHE_LINE_WID] mem_to_if_data;

MemCtrl mem_ctrl(
    .clk(clk_in),
    .rst(rst_in),
    .rdy(rdy_in),

    .rollback(rollback),

    .mem_din(mem_din),
    .mem_dout(mem_dout),
    .mem_a(mem_a),
    .mem_wr(mem_wr),

    .if_en(if_to_mem_en),
    .if_pc(if_to_mem_pc),
    .if_done(mem_to_if_done),
    .if_data(mem_to_if_data),

    .lsb_en(),
    .lsb_done()


);

IFetch(
    .clk,
    .rst,
    .rdy,

    .rollback,

    .rs_full,
    .lsb_full,
    .rob_full,

    .mem_en,
    .mem_pc,
    .mem_done,
    .mem_data,

    // now
    .inst_done,
    .inst,
    .inst_pc,
    .inst_pre_j,

    // when RoB commit
    .br_pre,
    .br_pre_j, // is jump
    .br_pre_pc,
    .br_res_pc
)

Decoder decoder(
    .clk(clk_in),
    .rst(rst_in),
    .rdy(rdy_in),

    .rollback(rollback),

    // fetch from IFetch
    .inst_done,
    .inst,
    .inst_pc,
    .inst_pre_j,

    // issue
    .done,
    .rob_pos,
    .opcode,
    .funct3,
    .funct7,
    .rs1_rdy,
    .rs1_val,
    .rs1_rob_pos,
    .rs2_rdy,
    .rs2_val,
    .rs2_rob_pos,
    .imm,
    .rd,
    .pc,
    .pre_j,

    // query from RegFile
    .reg_rs1,
    .reg_rs1_rdy,
    .reg_rs1_val,
    .reg_rs1_rob_pos,
    .reg_rs2,
    .reg_rs2_rdy,
    .reg_rs2_val,
    .reg_rs2_rob_pos,

    .rs_en,
    .lsb_en,

    .is_ready
);

endmodule